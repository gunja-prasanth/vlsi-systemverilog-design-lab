`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 16.02.2026 20:37:04
// Design Name: 
// Module Name: fsm_binary
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module fsm_binary (
    input  logic clk,
    input  logic rst,
    input  logic start,
    output logic done
);

    typedef enum logic [1:0] {
        IDLE    = 2'b00,
        LOAD    = 2'b01,
        PROCESS = 2'b10,
        DONE    = 2'b11
    } state_t;

    state_t current_state, next_state;

    always_ff @(posedge clk or posedge rst) begin
        if (rst)
            current_state <= IDLE;
        else
            current_state <= next_state;
    end

    always_comb begin
        next_state = current_state;
        done = 0;

        case (current_state)
            IDLE:    if (start) next_state = LOAD;
            LOAD:    next_state = PROCESS;
            PROCESS: next_state = DONE;
            DONE: begin
                done = 1;
                next_state = IDLE;
            end
        endcase
    end

endmodule
